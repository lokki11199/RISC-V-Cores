module adder (input  signed [31:0] a, //���� �� ��������� ���, ������������� wire? - ��
              input  signed [31:0] b,
              output signed [31:0] c
              );
              
assign c = a + b; //����������� ������������ - ������ �������������� ������
//� ��� ����� � ��� ����, ����� ������������ "signed"? - ��� ��������
//������������ �������� - ������������, �� �������, ��� ������� ��� ��������
              
endmodule